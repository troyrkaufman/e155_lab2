module hi()

endmodule